typedef virtual uart_if uart_vif;